library verilog;
use verilog.vl_types.all;
entity step_2_vlg_check_tst is
    port(
        F_POS           : in     vl_logic;
        F_SOP           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end step_2_vlg_check_tst;
