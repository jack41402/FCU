module step2(SW, KEY, HEX3, HEX2);
	input [9:2] SW;
	input [1:0] KEY;
	output reg[0:6] HEX3, HEX2;
	
	always @(SW, KEY) begin
		if (KEY[1]==0)
			case(SW[9:6])
				4'b0000: HEX3 = 7'b0000001;	// 0
				4'b0001: HEX3 = 7'b1001111;	// 1
				4'b0010: HEX3 = 7'b0010010;	// 2
				4'b0011: HEX3 = 7'b0000110;	// 3
				4'b0100: HEX3 = 7'b1001100;	// 4
				4'b0101: HEX3 = 7'b0100100;	// 5
				4'b0110: HEX3 = 7'b0100000;	// 6
				4'b0111: HEX3 = 7'b0001101;	// 7
				4'b1000: HEX3 = 7'b0000000;	// 8
				4'b1001: HEX3 = 7'b0000100;	// 9
				4'b1010: HEX3 = 7'b0001000;	// A
				4'b1011: HEX3 = 7'b1100000;	// B
				4'b1100: HEX3 = 7'b0110001;	// C
				4'b1101: HEX3 = 7'b1000010;	// D
				4'b1110: HEX3 = 7'b0110000;	// E
				4'b1111: HEX3 = 7'b0111000;	// F
				default: HEX3 = 7'b1111111; 	// default
			endcase
		else
			HEX3 = 7'b1111111;
		if (KEY[0]==0)
			case(SW[5:2])
				4'b0000: HEX2 = 7'b0000001;	// 0
				4'b0001: HEX2 = 7'b1001111;	// 1
				4'b0010: HEX2 = 7'b0010010;	// 2
				4'b0011: HEX2 = 7'b0000110;	// 3
				4'b0100: HEX2 = 7'b1001100;	// 4
				4'b0101: HEX2 = 7'b0100100;	// 5
				4'b0110: HEX2 = 7'b0100000;	// 6
				4'b0111: HEX2 = 7'b0001101;	// 7
				4'b1000: HEX2 = 7'b0000000;	// 8
				4'b1001: HEX2 = 7'b0000100;	// 9
				4'b1010: HEX2 = 7'b0001000;	// A
				4'b1011: HEX2 = 7'b1100000;	// B
				4'b1100: HEX2 = 7'b0110001;	// C
				4'b1101: HEX2 = 7'b1000010;	// D
				4'b1110: HEX2 = 7'b0110000;	// E
				4'b1111: HEX2 = 7'b0111000;	// F
				default: HEX2 = 7'b1111111; 	// default
			endcase
		else
			HEX2 = 7'b1111111;
	end
	
endmodule