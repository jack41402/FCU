library verilog;
use verilog.vl_types.all;
entity step1_vlg_vec_tst is
end step1_vlg_vec_tst;
