library verilog;
use verilog.vl_types.all;
entity step_2_vlg_vec_tst is
end step_2_vlg_vec_tst;
