module step1(v, d0, d1);
	input [3:0] v;
	output reg[0:6] d0, d1;
	
	always @(v) begin
		case(v)
			4'b0000, 4'b1010: d0 = 7'b0000001;	// 0
			4'b0001, 4'b1011: d0 = 7'b1001111;	// 1
			4'b0010, 4'b1100: d0 = 7'b0010010;	// 2
			4'b0011, 4'b1101: d0 = 7'b0000110;	// 3
			4'b0100, 4'b1110: d0 = 7'b1001100;	// 4
			4'b0101, 4'b1111: d0 = 7'b0100100;	// 5
			4'b0110			 : d0 = 7'b0100000;	// 6
			4'b0111			 : d0 = 7'b0001101;	// 7
			4'b1000			 : d0 = 7'b0000000;	// 8
			4'b1001			 : d0 = 7'b0000100;	// 9
			default			 : d0 = 7'b1111111;	// default
		endcase
		case(v)
			4'b0000, 4'b0001, 4'b0010,
			4'b0011, 4'b0100, 4'b0101,
			4'b0110, 4'b0111, 4'b1000, 4'b1001: d1 = 7'b0000001;	// 0
			
			4'b1010, 4'b1011, 4'b1100,
			4'b1101, 4'b1110, 4'b1111			 : d1 = 7'b1001111;	// 1
			default			 						 : d1 = 7'b1111111;	// default
		endcase
	end
endmodule