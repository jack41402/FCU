library verilog;
use verilog.vl_types.all;
entity step_1_vlg_vec_tst is
end step_1_vlg_vec_tst;
